*mat_array.cir


*Row Voltage Sources
V1 RowC_1 0 -5.000000
V3 RowC_2 0 -5.000000


*Row Current Sources
I1 I_1 0 -0.000000
I3 I_3 0 -0.000000


*Row 'Ammeter' Resistances
R41 RowC_1 MemRRow4 0.000000001000
R42 RowC_2 MemRRow7 0.000000001000


*Memristor Resistances
R14 MemRRow4 MemRCol4 6666670.000000
R18 MemRRow8 MemRCol8 3333340.000000
R17 MemRRow7 MemRCol7 3333340.000000
R112 MemRRow12 MemRCol12 10.000000


*Line Row Resistances
R24 MemRRow4 MemRRow8 10.000000
R28 MemRRow8 MemRRow13 10.000000
R27 MemRRow7 MemRRow12 10.000000
R212 MemRRow12 MemRRow18 10.000000


*Line Column Resistances
R34 MemRCol4 MemRCol7 10.000000
R38 MemRCol8 MemRCol12 10.000000
R37 MemRCol7 MemRCol11 10.000000
R312 MemRCol12 MemRCol17 10.000000


*Column 'Ammeter' Resistances
R51 MemRCol11 ColC_1 0.000000001000
R52 MemRCol17 ColC_2 0.000000001000


*Column Voltage Sources
V2 ColC_1 0 0.000000
V5 ColC_2 0 0.000000


*Column Current Sources
I2 I_2 0 -0.000000
I5 I_5 0 -0.000000


*Spice Directives
.op
*.backanno
.end
