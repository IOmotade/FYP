*mat_array.cir


*Voltage Sources
V1 V_1 0 5.000000
V2 V_2 0 5.000000
V3 V_3 0 5.000000


*Row 'Ammeter' Resistances
R41 V_1 MemRRow11 0.000000001000
R42 V_2 MemRRow21 0.000000001000
R43 V_3 MemRRow31 0.000000001000


*Memristor Resistances
R14 MemRRow4 MemRCol4 10000.000000
R18 MemRRow8 MemRCol8 10000.000000
R113 MemRRow13 MemRCol13 10000.000000
R17 MemRRow7 MemRCol7 10000.000000
R112 MemRRow12 MemRCol12 10000.000000
R118 MemRRow18 MemRCol18 10000.000000
R111 MemRRow11 MemRCol11 10000.000000
R117 MemRRow17 MemRCol17 10000.000000
R124 MemRRow24 MemRCol24 10000.000000


*Line Row Resistances
R24 MemRRow4 MemRRow8 1000.000000
R28 MemRRow8 MemRRow13 1000.000000
R213 MemRRow13 MemRRow19 1000.000000
R27 MemRRow7 MemRRow12 1000.000000
R212 MemRRow12 MemRRow18 1000.000000
R218 MemRRow18 MemRRow25 1000.000000
R211 MemRRow11 MemRRow17 1000.000000
R217 MemRRow17 MemRRow24 1000.000000
R224 MemRRow24 MemRRow32 1000.000000


*Line Column Resistances
R34 MemRCol4 MemRCol7 1000.000000
R38 MemRCol8 MemRCol12 1000.000000
R313 MemRCol13 MemRCol18 1000.000000
R37 MemRCol7 MemRCol11 1000.000000
R312 MemRCol12 MemRCol17 1000.000000
R318 MemRCol18 MemRCol24 1000.000000
R311 MemRCol11 MemRCol16 1000.000000
R317 MemRCol17 MemRCol23 1000.000000
R324 MemRCol24 MemRCol31 1000.000000


*Column 'Ammeter' Resistances
R51 MemRCol16 0 0.000000001000
R52 MemRCol23 0 0.000000001000
R53 MemRCol31 0 0.000000001000


*Spice Directives
.op
*.backanno
.end
